.SUBCKT ASYNC_DFFHx1_ASAP7_75t_R CLK D QN RESET SET VDD VSS
MMMMMMMMMMM43 1 SET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMM24 QN SH VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMM29 SS SH VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMM23 clkb clkn VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMM20 clkn CLK VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMM44 SS RESET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMM34 SH clkn 1 VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMM48 net020 RESET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMM12 MS clkb SH VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMM33 1 SS VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMM9 MH clkb net020 VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMM8 net020 MS VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMM6 MS MH VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMM5 pd1 D VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMM4 MH clkn pd1 VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMM47 MS SET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMM25 QN SH VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMM28 SS SH net076 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMM22 clkb clkn VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMM45 net076 RESET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMM46 net079 SET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMM21 clkn CLK VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMM37 2 SS net077 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMM35 SH clkb 2 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMM49 net078 RESET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMM13 MS clkn SH VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMM11 net051 MS net078 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMM10 MH clkn net051 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMM7 MS MH net079 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMM42 net077 SET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMM1 MH clkb pu1 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMM3 pu1 D VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMM43 pd3 SET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMM24 QN SH VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMM29 SS SH VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMM23 clkb clkn VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMM20 clkn CLK VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMM44 SS RESET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMM34 SH clkn pd3 VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMM48 net020 RESET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMM12 MS clkb SH VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMM33 3 SS VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMM9 MH clkb 7 VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMM8 7 MS VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMM6 MS MH VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMM5 13 D VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMM4 MH clkn 13 VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMM47 MS SET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMM25 QN SH VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMM28 SS SH net076 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMM22 clkb clkn VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMM45 net076 RESET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMM46 net079 SET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMM21 clkn CLK VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMM37 2 SS net077 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMM35 SH clkb 12 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMM49 net078 RESET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMM13 MS clkn SH VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMM11 net051 MS net078 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMM10 MH clkn net051 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMM7 MS MH net079 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMM42 net077 SET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMM1 MH clkb pu1 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMM3 pu1 D VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMM43 3 SET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMM24 QN SH VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMM29 SS SH VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMM23 clkb clkn VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMM20 clkn CLK VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMM44 SS RESET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMM34 SH clkn 3 VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMM48 7 RESET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMM12 MS clkb SH VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMM33 14 SS VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMM9 MH clkb 4 VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMM8 4 MS VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMM6 MS MH VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMM5 13 D VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMM4 MH clkn 13 VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMM47 MS SET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMM25 QN SH VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMM28 SS SH net076 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMM22 clkb clkn VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMM45 8 RESET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMM46 net079 SET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMM21 clkn CLK VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMM37 pd2 SS 5 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMM35 SH clkb 15 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMM49 net078 RESET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMM13 MS clkn SH VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMM11 net051 MS net078 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMM10 MH clkn net051 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMM7 MS MH net079 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMM42 5 SET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMM1 MH clkb pu1 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMM3 pu1 D VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMM43 14 SET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMM24 QN SH VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMM29 SS SH VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMM23 clkb clkn VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMM20 clkn CLK VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMM44 SS RESET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMM34 SH clkn 14 VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMM48 4 RESET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMM12 MS clkb SH VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMM33 16 SS VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMM9 MH clkb 4 VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMM8 6 MS VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMM6 MS MH VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMM5 pd1 D VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMM4 MH clkn pd1 VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMM47 MS SET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMM25 QN SH VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMM28 SS SH 8 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMM22 clkb clkn VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMM45 8 RESET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMM46 net079 SET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMM21 clkn CLK VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMM37 15 SS 5 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMM35 SH clkb 15 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMM49 net078 RESET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMM13 MS clkn SH VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMM11 net051 MS net078 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMM10 MH clkn net051 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMM7 MS MH net079 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMM42 net077 SET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMM1 MH clkb pu1 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMM3 pu1 D VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMM43 16 SET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMM24 QN SH VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMM29 SS SH VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMM23 clkb clkn VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMM20 clkn CLK VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMM44 SS RESET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMM34 SH clkn 16 VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMM48 6 RESET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMM12 MS clkb SH VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMM33 pd3 SS VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMM9 MH clkb 6 VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMM8 net020 MS VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMM6 MS MH VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMM5 pd1 D VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMM4 MH clkn pd1 VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMM47 MS SET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMM25 QN SH VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMM28 SS SH net076 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMM22 clkb clkn VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMM45 net076 RESET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMM46 net079 SET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMM21 clkn CLK VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMM37 pd2 SS net077 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMM35 SH clkb pd2 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMM49 net078 RESET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMM13 MS clkn SH VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMM11 9 MS net078 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMM10 MH clkn 9 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMM7 MS MH net079 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMM42 net077 SET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMM1 MH clkb pu1 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMM3 pu1 D VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMMM43 pd3 SET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMMM24 QN SH VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMMM29 SS SH VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMMM23 clkb clkn VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMMM20 clkn CLK VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMMM44 SS RESET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMMM34 SH clkn pd3 VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMMM48 net020 RESET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMMM12 MS clkb SH VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMMM33 pd3 SS VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMMM9 MH clkb net020 VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMMM8 net020 MS VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMMM6 MS MH VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMMM5 pd1 D VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMMM4 MH clkn pd1 VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMMM47 MS SET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMMM25 QN SH VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMMM28 SS SH 10 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMMM22 clkb clkn VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMMM45 10 RESET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMMM46 net079 SET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMMM21 clkn CLK VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMMM37 pd2 SS net077 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMMM35 SH clkb 12 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMMM49 net078 RESET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMMM13 MS clkn SH VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMMM11 9 MS net078 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMMM10 MH clkn net051 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMMM7 MS MH net079 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMMM42 net077 SET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMMM1 MH clkb pu1 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMMM3 pu1 D VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMMMM43 11 SET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMMMM24 QN SH VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMMMM29 SS SH VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMMMM23 clkb clkn VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMMMM20 clkn CLK VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMMMM44 SS RESET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMMMM34 SH clkn 11 VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMMMM48 net020 RESET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMMMM12 MS clkb SH VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMMMM33 11 SS VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMMMM9 MH clkb net020 VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMMMM8 net020 MS VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMMMM6 MS MH VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMMMM5 pd1 D VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMMMM4 MH clkn pd1 VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMMMM47 MS SET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMMMMMMMMMMMMMMMMMMM25 QN SH VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMMMM28 SS SH 10 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMMMM22 clkb clkn VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMMMM45 net076 RESET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMMMM46 net079 SET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMMMM21 clkn CLK VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMMMM37 12 SS net077 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMMMM35 SH clkb 12 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMMMM49 net078 RESET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMMMM13 MS clkn SH VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMMMM11 net051 MS net078 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMMMM10 MH clkn net051 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMMMM7 MS MH net079 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMMMM42 net077 SET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMMMM1 MH clkb pu1 VDD pmos_rvt w=162.0n l=20n nfin=6
MMMMMMMMMMMMMMMMMMMM3 pu1 D VDD VDD pmos_rvt w=162.0n l=20n nfin=6
.ENDS